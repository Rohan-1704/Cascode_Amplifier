magic
tech scmos
timestamp 1699373897
<< nwell >>
rect -28 -4 66 63
<< ntransistor >>
rect 13 -37 18 -17
rect 13 -77 18 -57
<< ptransistor >>
rect -4 6 0 50
rect 41 6 45 50
<< ndiffusion >>
rect -1 -28 13 -17
rect -1 -34 1 -28
rect 8 -34 13 -28
rect -1 -37 13 -34
rect 18 -22 31 -17
rect 18 -29 23 -22
rect 29 -29 31 -22
rect 18 -37 31 -29
rect -1 -64 13 -57
rect -1 -70 1 -64
rect 8 -70 13 -64
rect -1 -77 13 -70
rect 18 -65 31 -57
rect 18 -72 21 -65
rect 28 -72 31 -65
rect 18 -77 31 -72
<< pdiffusion >>
rect -11 47 -4 50
rect -11 42 -10 47
rect -6 42 -4 47
rect -11 6 -4 42
rect 0 47 7 50
rect 0 42 2 47
rect 6 42 7 47
rect 0 6 7 42
rect 34 47 41 50
rect 34 42 35 47
rect 39 42 41 47
rect 34 6 41 42
rect 45 14 55 50
rect 45 9 49 14
rect 53 9 55 14
rect 45 6 55 9
<< ndcontact >>
rect 1 -34 8 -28
rect 23 -29 29 -22
rect 1 -70 8 -64
rect 21 -72 28 -65
<< pdcontact >>
rect -10 42 -6 47
rect 2 42 6 47
rect 35 42 39 47
rect 49 9 53 14
<< psubstratepcontact >>
rect -13 -99 -8 -94
rect 1 -99 6 -94
rect 14 -99 19 -94
rect 29 -99 34 -94
rect 41 -99 46 -94
<< nsubstratencontact >>
rect -15 56 -10 60
rect 4 56 9 60
rect 18 56 23 60
rect 32 56 37 60
rect 45 56 50 60
<< polycontact >>
rect -8 0 -4 4
rect 37 0 41 4
rect 18 -44 23 -39
rect 9 -84 13 -79
<< polypplus >>
rect -4 50 0 53
rect 41 50 45 53
rect -4 0 0 6
rect 41 0 45 6
rect 13 -41 18 -40
<< polynplus >>
rect 13 -17 18 -12
rect 13 -40 18 -37
rect 13 -44 18 -41
rect 13 -57 18 -52
rect 13 -84 18 -77
<< metal1 >>
rect -21 60 56 61
rect -21 56 -15 60
rect -10 56 4 60
rect 9 56 18 60
rect 23 56 32 60
rect 37 56 45 60
rect 50 56 56 60
rect -10 47 -6 56
rect 6 42 35 47
rect 39 42 40 47
rect 48 14 54 17
rect 48 9 49 14
rect 53 9 54 14
rect -19 4 0 6
rect -19 0 -8 4
rect -4 0 0 4
rect 26 4 45 6
rect 26 0 37 4
rect 41 0 45 4
rect 48 -22 54 9
rect 29 -29 54 -22
rect 1 -64 8 -34
rect 13 -44 18 -39
rect 23 -44 29 -39
rect 2 -84 9 -79
rect 13 -84 18 -79
rect 21 -92 28 -72
rect -16 -94 53 -92
rect -16 -99 -13 -94
rect -8 -99 1 -94
rect 6 -99 14 -94
rect 19 -99 29 -94
rect 34 -99 41 -94
rect 46 -99 53 -94
rect -16 -100 53 -99
<< labels >>
rlabel metal1 24 58 24 58 5 VDD
rlabel space 30 -42 30 -42 1 Vbias3
rlabel metal1 26 3 26 3 1 Vbias2
rlabel nwell -20 3 -20 3 1 Vbias1
rlabel metal1 5 -82 5 -82 1 Vin
rlabel metal1 10 -97 10 -97 1 GND
<< end >>
